`default_nettype none

module mod_WarpScheduler();
    // Placeholder
endmodule
